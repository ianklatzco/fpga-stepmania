
module audio (
	clk_clk,
	reset_reset_n,
	pll_clk_out_18mhz_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		pll_clk_out_18mhz_clk;
endmodule
