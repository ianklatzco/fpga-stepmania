/*module(

);*/