Dashiell                                              D a s h i e l l       	 M S   G o t h i c          � �              � �                           