module audio_loop (
	input  logic Clk,
	input  logic reset,
	output logic [15:0] audio_data
);

logic [15:0] mem [0:999];

// $readmemb("piano.wav",mem); // only works in testbenching, which we don't care about

int counter = 0;
// playback of ROM
always_ff @(posedge Clk or posedge reset)
begin
	if(reset) begin
		counter <= 0;
	end else begin
		if (counter >= 1000) begin
			audio_data <= mem[0];
			counter <= 0;
		end else begin
		 	audio_data <= mem[counter];
			counter <= counter + 1;
		end
	end
end

// loading BRAM with a ROM containing a simple alternating pulse
// copied from lab6 and modifed to our needs
always_ff @ (posedge Clk or posedge reset)
begin
	if(reset)
	begin
// mem[0] <= 16'hf3ff;
// mem[1] <= 16'h0000;
// mem[2] <= 16'hf0ff;
// mem[3] <= 16'h0000;
// mem[4] <= 16'hfbff;
// mem[5] <= 16'hf1ff;
// mem[6] <= 16'hffff;
// mem[7] <= 16'hffff;
// mem[8] <= 16'hf9ff;
// mem[9] <= 16'hf7ff;
// mem[10] <= 16'hf7ff;
// mem[11] <= 16'hf3ff;
// mem[12] <= 16'hffff;
// mem[13] <= 16'hfdff;
// mem[14] <= 16'hfbff;
// mem[15] <= 16'hf9ff;
// mem[16] <= 16'hfbff;
// mem[17] <= 16'hf9ff;
// mem[18] <= 16'hffff;
// mem[19] <= 16'hfbff;
// mem[20] <= 16'hfdff;
// mem[21] <= 16'hf9ff;
// mem[22] <= 16'hfdff;
// mem[23] <= 16'hf2ff;
// mem[24] <= 16'hffff;
// mem[25] <= 16'hffff;
// mem[26] <= 16'hfbff;
// mem[27] <= 16'hfbff;
// mem[28] <= 16'h0200;
// mem[29] <= 16'hf5ff;
// mem[30] <= 16'hfbff;
// mem[31] <= 16'hffff;
// mem[32] <= 16'hfbff;
// mem[33] <= 16'hf9ff;
// mem[34] <= 16'hf5ff;
// mem[35] <= 16'h0000;
// mem[36] <= 16'hf9ff;
// mem[37] <= 16'hfdff;
// mem[38] <= 16'hf9ff;
// mem[39] <= 16'hf9ff;
// mem[40] <= 16'hf9ff;
// mem[41] <= 16'h0000;
// mem[42] <= 16'hf7ff;
// mem[43] <= 16'hf5ff;
// mem[44] <= 16'hffff;
// mem[45] <= 16'hf2ff;
// mem[46] <= 16'h0000;
// mem[47] <= 16'hffff;
// mem[48] <= 16'hfbff;
// mem[49] <= 16'hffff;
// mem[50] <= 16'hf5ff;
// mem[51] <= 16'hffff;
// mem[52] <= 16'hf3ff;
// mem[53] <= 16'h0300;
// mem[54] <= 16'hfbff;
// mem[55] <= 16'hf5ff;
// mem[56] <= 16'hffff;
// mem[57] <= 16'hf9ff;
// mem[58] <= 16'hfbff;
// mem[59] <= 16'hf7ff;
// mem[60] <= 16'hffff;
// mem[61] <= 16'hfbff;
// mem[62] <= 16'hfdff;
// mem[63] <= 16'hffff;
// mem[64] <= 16'hf2ff;
// mem[65] <= 16'hfdff;
// mem[66] <= 16'hfbff;
// mem[67] <= 16'hf9ff;
// mem[68] <= 16'hf7ff;
// mem[69] <= 16'hf9ff;
// mem[70] <= 16'hf7ff;
// mem[71] <= 16'hfdff;
// mem[72] <= 16'hfdff;
// mem[73] <= 16'hf9ff;
// mem[74] <= 16'hffff;
// mem[75] <= 16'hfbff;
// mem[76] <= 16'hffff;
// mem[77] <= 16'hf7ff;
// mem[78] <= 16'hfdff;
// mem[79] <= 16'hf9ff;
// mem[80] <= 16'hf0ff;
// mem[81] <= 16'h0700;
// mem[82] <= 16'hf9ff;
// mem[83] <= 16'hfbff;
// mem[84] <= 16'hfbff;
// mem[85] <= 16'hfdff;
// mem[86] <= 16'hf9ff;
// mem[87] <= 16'hf9ff;
// mem[88] <= 16'hf9ff;
// mem[89] <= 16'h0300;
// mem[90] <= 16'hfdff;
// mem[91] <= 16'hfdff;
// mem[92] <= 16'hfdff;
// mem[93] <= 16'hffff;
// mem[94] <= 16'hffff;
// mem[95] <= 16'hf9ff;
// mem[96] <= 16'hfbff;
// mem[97] <= 16'h0200;
// mem[98] <= 16'hffff;
// mem[99] <= 16'hffff;
// mem[100] <= 16'h0000;
// mem[101] <= 16'h0200;
// mem[102] <= 16'hffff;
// mem[103] <= 16'hfdff;
// mem[104] <= 16'h0400;
// mem[105] <= 16'hfdff;
// mem[106] <= 16'hfdff;
// mem[107] <= 16'h0000;
// mem[108] <= 16'hfbff;
// mem[109] <= 16'hfdff;
// mem[110] <= 16'hfdff;
// mem[111] <= 16'h0200;
// mem[112] <= 16'hf2ff;
// mem[113] <= 16'h0500;
// mem[114] <= 16'hf7ff;
// mem[115] <= 16'h0700;
// mem[116] <= 16'hf9ff;
// mem[117] <= 16'hf9ff;
// mem[118] <= 16'h0700;
// mem[119] <= 16'hf9ff;
// mem[120] <= 16'h0200;
// mem[121] <= 16'h0200;
// mem[122] <= 16'hfbff;
// mem[123] <= 16'hfbff;
// mem[124] <= 16'h0700;
// mem[125] <= 16'hfdff;
// mem[126] <= 16'h0300;
// mem[127] <= 16'hf9ff;
// mem[128] <= 16'h0400;
// mem[129] <= 16'hfdff;
// mem[130] <= 16'hfdff;
// mem[131] <= 16'h0900;
// mem[132] <= 16'hf7ff;
// mem[133] <= 16'h0500;
// mem[134] <= 16'h0300;
// mem[135] <= 16'hfdff;
// mem[136] <= 16'h0200;
// mem[137] <= 16'hfdff;
// mem[138] <= 16'hfdff;
// mem[139] <= 16'h0400;
// mem[140] <= 16'hffff;
// mem[141] <= 16'h0500;
// mem[142] <= 16'hfbff;
// mem[143] <= 16'hfdff;
// mem[144] <= 16'h0900;
// mem[145] <= 16'h0200;
// mem[146] <= 16'h0200;
// mem[147] <= 16'hffff;
// mem[148] <= 16'h0200;
// mem[149] <= 16'h0300;
// mem[150] <= 16'h0000;
// mem[151] <= 16'h0d00;
// mem[152] <= 16'hfdff;
// mem[153] <= 16'hfdff;
// mem[154] <= 16'h0000;
// mem[155] <= 16'h0500;
// mem[156] <= 16'h0200;
// mem[157] <= 16'h0500;
// mem[158] <= 16'hfdff;
// mem[159] <= 16'h0400;
// mem[160] <= 16'h0900;
// mem[161] <= 16'h0500;
// mem[162] <= 16'h0500;
// mem[163] <= 16'h0700;
// mem[164] <= 16'h0000;
// mem[165] <= 16'h0000;
// mem[166] <= 16'h0f00;
// mem[167] <= 16'hfdff;
// mem[168] <= 16'h0900;
// mem[169] <= 16'h0300;
// mem[170] <= 16'h0700;
// mem[171] <= 16'h0900;
// mem[172] <= 16'h0700;
// mem[173] <= 16'hfdff;
// mem[174] <= 16'h0700;
// mem[175] <= 16'h0700;
// mem[176] <= 16'h0000;
// mem[177] <= 16'h0000;
// mem[178] <= 16'h0500;
// mem[179] <= 16'h0500;
// mem[180] <= 16'h0500;
// mem[181] <= 16'h0500;
// mem[182] <= 16'h0000;
// mem[183] <= 16'h0900;
// mem[184] <= 16'h0900;
// mem[185] <= 16'h0500;
// mem[186] <= 16'h0400;
// mem[187] <= 16'h0900;
// mem[188] <= 16'h0200;
// mem[189] <= 16'h0500;
// mem[190] <= 16'h0500;
// mem[191] <= 16'h0200;
// mem[192] <= 16'h0b00;
// mem[193] <= 16'h0500;
// mem[194] <= 16'h0500;
// mem[195] <= 16'h0200;
// mem[196] <= 16'h0d00;
// mem[197] <= 16'h0200;
// mem[198] <= 16'h0200;
// mem[199] <= 16'h0b00;
// mem[200] <= 16'h0700;
// mem[201] <= 16'hffff;
// mem[202] <= 16'h0b00;
// mem[203] <= 16'h0b00;
// mem[204] <= 16'h0500;
// mem[205] <= 16'h0200;
// mem[206] <= 16'h0200;
// mem[207] <= 16'h0700;
// mem[208] <= 16'hfdff;
// mem[209] <= 16'h0b00;
// mem[210] <= 16'h0700;
// mem[211] <= 16'hffff;
// mem[212] <= 16'h0500;
// mem[213] <= 16'h0700;
// mem[214] <= 16'h0400;
// mem[215] <= 16'h0500;
// mem[216] <= 16'h0500;
// mem[217] <= 16'hffff;
// mem[218] <= 16'h0b00;
// mem[219] <= 16'h0400;
// mem[220] <= 16'h0400;
// mem[221] <= 16'h0000;
// mem[222] <= 16'h0400;
// mem[223] <= 16'h0200;
// mem[224] <= 16'h0400;
// mem[225] <= 16'h0200;
// mem[226] <= 16'h0200;
// mem[227] <= 16'h0300;
// mem[228] <= 16'hffff;
// mem[229] <= 16'h0500;
// mem[230] <= 16'h0300;
// mem[231] <= 16'hfbff;
// mem[232] <= 16'h0500;
// mem[233] <= 16'h0400;
// mem[234] <= 16'h0200;
// mem[235] <= 16'h0000;
// mem[236] <= 16'hfdff;
// mem[237] <= 16'h0300;
// mem[238] <= 16'hfbff;
// mem[239] <= 16'hffff;
// mem[240] <= 16'h0700;
// mem[241] <= 16'h0200;
// mem[242] <= 16'hfdff;
// mem[243] <= 16'h0500;
// mem[244] <= 16'h0400;
// mem[245] <= 16'h0200;
// mem[246] <= 16'h0300;
// mem[247] <= 16'hffff;
// mem[248] <= 16'h0600;
// mem[249] <= 16'h0200;
// mem[250] <= 16'h0300;
// mem[251] <= 16'hffff;
// mem[252] <= 16'h0200;
// mem[253] <= 16'hffff;
// mem[254] <= 16'hffff;
// mem[255] <= 16'h0000;
// mem[256] <= 16'hfcff;
// mem[257] <= 16'hf7ff;
// mem[258] <= 16'h0600;
// mem[259] <= 16'hffff;
// mem[260] <= 16'h0200;
// mem[261] <= 16'h0200;
// mem[262] <= 16'hfdff;
// mem[263] <= 16'hffff;
// mem[264] <= 16'hffff;
// mem[265] <= 16'h0400;
// mem[266] <= 16'hf9ff;
// mem[267] <= 16'h0000;
// mem[268] <= 16'h0300;
// mem[269] <= 16'h0000;
// mem[270] <= 16'h0300;
// mem[271] <= 16'h0200;
// mem[272] <= 16'h0000;
// mem[273] <= 16'hf9ff;
// mem[274] <= 16'hfdff;
// mem[275] <= 16'hffff;
// mem[276] <= 16'h0200;
// mem[277] <= 16'hffff;
// mem[278] <= 16'hf7ff;
// mem[279] <= 16'h0700;
// mem[280] <= 16'h0000;
// mem[281] <= 16'hffff;
// mem[282] <= 16'h0300;
// mem[283] <= 16'h0000;
// mem[284] <= 16'hffff;
// mem[285] <= 16'h0000;
// mem[286] <= 16'h0000;
// mem[287] <= 16'h0200;
// mem[288] <= 16'hf5ff;
// mem[289] <= 16'h0300;
// mem[290] <= 16'h0300;
// mem[291] <= 16'hffff;
// mem[292] <= 16'h0000;
// mem[293] <= 16'hffff;
// mem[294] <= 16'h0000;
// mem[295] <= 16'hfdff;
// mem[296] <= 16'hffff;
// mem[297] <= 16'hfbff;
// mem[298] <= 16'h0000;
// mem[299] <= 16'hfbff;
// mem[300] <= 16'hfdff;
// mem[301] <= 16'hf9ff;
// mem[302] <= 16'h0200;
// mem[303] <= 16'hfdff;
// mem[304] <= 16'hfdff;
// mem[305] <= 16'hffff;
// mem[306] <= 16'hf7ff;
// mem[307] <= 16'h0500;
// mem[308] <= 16'hf9ff;
// mem[309] <= 16'hffff;
// mem[310] <= 16'hfdff;
// mem[311] <= 16'hfbff;
// mem[312] <= 16'hfbff;
// mem[313] <= 16'hffff;
// mem[314] <= 16'hf9ff;
// mem[315] <= 16'h0000;
// mem[316] <= 16'hf5ff;
// mem[317] <= 16'hffff;
// mem[318] <= 16'h0200;
// mem[319] <= 16'hffff;
// mem[320] <= 16'hfdff;
// mem[321] <= 16'hfbff;
// mem[322] <= 16'hfbff;
// mem[323] <= 16'h0000;
// mem[324] <= 16'hfdff;
// mem[325] <= 16'hfdff;
// mem[326] <= 16'hffff;
// mem[327] <= 16'hfdff;
// mem[328] <= 16'hffff;
// mem[329] <= 16'hfdff;
// mem[330] <= 16'hffff;
// mem[331] <= 16'hfdff;
// mem[332] <= 16'hf3ff;
// mem[333] <= 16'h0200;
// mem[334] <= 16'hfdff;
// mem[335] <= 16'h0400;
// mem[336] <= 16'hf7ff;
// mem[337] <= 16'hfdff;
// mem[338] <= 16'hffff;
// mem[339] <= 16'hffff;
// mem[340] <= 16'hfbff;
// mem[341] <= 16'hffff;
// mem[342] <= 16'hffff;
// mem[343] <= 16'hffff;
// mem[344] <= 16'hf1ff;
// mem[345] <= 16'h0200;
// mem[346] <= 16'h0000;
// mem[347] <= 16'hf9ff;
// mem[348] <= 16'hfbff;
// mem[349] <= 16'hf9ff;
// mem[350] <= 16'h0000;
// mem[351] <= 16'h0200;
// mem[352] <= 16'h0000;
// mem[353] <= 16'hf7ff;
// mem[354] <= 16'hfbff;
// mem[355] <= 16'h0300;
// mem[356] <= 16'hfbff;
// mem[357] <= 16'hffff;
// mem[358] <= 16'hfdff;
// mem[359] <= 16'hfbff;
// mem[360] <= 16'hf3ff;
// mem[361] <= 16'h0400;
// mem[362] <= 16'hfdff;
// mem[363] <= 16'hffff;
// mem[364] <= 16'hfbff;
// mem[365] <= 16'hfdff;
// mem[366] <= 16'hf9ff;
// mem[367] <= 16'hfdff;
// mem[368] <= 16'h0000;
// mem[369] <= 16'hfbff;
// mem[370] <= 16'hf5ff;
// mem[371] <= 16'hffff;
// mem[372] <= 16'hf7ff;
// mem[373] <= 16'h0000;
// mem[374] <= 16'hf5ff;
// mem[375] <= 16'h0300;
// mem[376] <= 16'hf9ff;
// mem[377] <= 16'hfbff;
// mem[378] <= 16'hffff;
// mem[379] <= 16'hfbff;
// mem[380] <= 16'h0000;
// mem[381] <= 16'hfbff;
// mem[382] <= 16'hfbff;
// mem[383] <= 16'hffff;
// mem[384] <= 16'hfeff;
// mem[385] <= 16'hfbff;
// mem[386] <= 16'hfdff;
// mem[387] <= 16'hfdff;
// mem[388] <= 16'hfdff;
// mem[389] <= 16'hfdff;
// mem[390] <= 16'hfdff;
// mem[391] <= 16'hfdff;
// mem[392] <= 16'hf9ff;
// mem[393] <= 16'hffff;
// mem[394] <= 16'hfbff;
// mem[395] <= 16'hf9ff;
// mem[396] <= 16'h0200;
// mem[397] <= 16'hfdff;
// mem[398] <= 16'hfdff;
// mem[399] <= 16'hfdff;
// mem[400] <= 16'hfdff;
// mem[401] <= 16'hf9ff;
// mem[402] <= 16'hfdff;
// mem[403] <= 16'hfdff;
// mem[404] <= 16'hfbff;
// mem[405] <= 16'hf9ff;
// mem[406] <= 16'hfdff;
// mem[407] <= 16'hfdff;
// mem[408] <= 16'hfdff;
// mem[409] <= 16'hfbff;
// mem[410] <= 16'hfdff;
// mem[411] <= 16'hfdff;
// mem[412] <= 16'hf5ff;
// mem[413] <= 16'h0000;
// mem[414] <= 16'hffff;
// mem[415] <= 16'hf9ff;
// mem[416] <= 16'h0200;
// mem[417] <= 16'hf3ff;
// mem[418] <= 16'hf9ff;
// mem[419] <= 16'hfdff;
// mem[420] <= 16'hfdff;
// mem[421] <= 16'hfdff;
// mem[422] <= 16'hfdff;
// mem[423] <= 16'hfdff;
// mem[424] <= 16'hfbff;
// mem[425] <= 16'hfbff;
// mem[426] <= 16'hfdff;
// mem[427] <= 16'hfdff;
// mem[428] <= 16'hfbff;
// mem[429] <= 16'hfdff;
// mem[430] <= 16'h0000;
// mem[431] <= 16'hf1ff;
// mem[432] <= 16'hf9ff;
// mem[433] <= 16'hfdff;
// mem[434] <= 16'hfbff;
// mem[435] <= 16'hfbff;
// mem[436] <= 16'hf7ff;
// mem[437] <= 16'hfbff;
// mem[438] <= 16'hffff;
// mem[439] <= 16'hf1ff;
// mem[440] <= 16'hfbff;
// mem[441] <= 16'hf9ff;
// mem[442] <= 16'hf9ff;
// mem[443] <= 16'hffff;
// mem[444] <= 16'hfdff;
// mem[445] <= 16'hf7ff;
// mem[446] <= 16'hfbff;
// mem[447] <= 16'hfbff;
// mem[448] <= 16'hf5ff;
// mem[449] <= 16'h0000;
// mem[450] <= 16'hf5ff;
// mem[451] <= 16'hf5ff;
// mem[452] <= 16'hffff;
// mem[453] <= 16'hf9ff;
// mem[454] <= 16'hfbff;
// mem[455] <= 16'hfbff;
// mem[456] <= 16'hfdff;
// mem[457] <= 16'hf9ff;
// mem[458] <= 16'hfbff;
// mem[459] <= 16'hf9ff;
// mem[460] <= 16'hfbff;
// mem[461] <= 16'hf1ff;
// mem[462] <= 16'hffff;
// mem[463] <= 16'hf7ff;
// mem[464] <= 16'hf7ff;
// mem[465] <= 16'hfbff;
// mem[466] <= 16'hfbff;
// mem[467] <= 16'hf3ff;
// mem[468] <= 16'hf9ff;
// mem[469] <= 16'hfdff;
// mem[470] <= 16'hf5ff;
// mem[471] <= 16'hf7ff;
// mem[472] <= 16'hffff;
// mem[473] <= 16'hf7ff;
// mem[474] <= 16'hfbff;
// mem[475] <= 16'hf7ff;
// mem[476] <= 16'hffff;
// mem[477] <= 16'hf5ff;
// mem[478] <= 16'hf5ff;
// mem[479] <= 16'h0000;
// mem[480] <= 16'hf5ff;
// mem[481] <= 16'hfdff;
// mem[482] <= 16'hf5ff;
// mem[483] <= 16'hffff;
// mem[484] <= 16'hffff;
// mem[485] <= 16'hf9ff;
// mem[486] <= 16'hf9ff;
// mem[487] <= 16'hffff;
// mem[488] <= 16'hfdff;
// mem[489] <= 16'hfbff;
// mem[490] <= 16'hffff;
// mem[491] <= 16'hf5ff;
// mem[492] <= 16'hfeff;
// mem[493] <= 16'h0000;
// mem[494] <= 16'hf3ff;
// mem[495] <= 16'hfdff;
// mem[496] <= 16'hfdff;
// mem[497] <= 16'hf5ff;
// mem[498] <= 16'hfbff;
// mem[499] <= 16'hf5ff;
// mem[500] <= 16'hfbff;
// mem[501] <= 16'hfdff;
// mem[502] <= 16'hfbff;
// mem[503] <= 16'hf9ff;
// mem[504] <= 16'hfdff;
// mem[505] <= 16'hf7ff;
// mem[506] <= 16'hffff;
// mem[507] <= 16'hf5ff;
// mem[508] <= 16'hfeff;
// mem[509] <= 16'h0200;
// mem[510] <= 16'hfeff;
// mem[511] <= 16'hf9ff;
// mem[512] <= 16'hfdff;
// mem[513] <= 16'hf5ff;
// mem[514] <= 16'h0000;
// mem[515] <= 16'hf9ff;
// mem[516] <= 16'hfbff;
// mem[517] <= 16'hffff;
// mem[518] <= 16'h0000;
// mem[519] <= 16'hffff;
// mem[520] <= 16'hffff;
// mem[521] <= 16'hfbff;
// mem[522] <= 16'hfdff;
// mem[523] <= 16'hfbff;
// mem[524] <= 16'hf7ff;
// mem[525] <= 16'h0500;
// mem[526] <= 16'hfdff;
// mem[527] <= 16'h0200;
// mem[528] <= 16'hffff;
// mem[529] <= 16'hf9ff;
// mem[530] <= 16'h0300;
// mem[531] <= 16'h0000;
// mem[532] <= 16'hfbff;
// mem[533] <= 16'hffff;
// mem[534] <= 16'h0500;
// mem[535] <= 16'hfdff;
// mem[536] <= 16'h0400;
// mem[537] <= 16'hffff;
// mem[538] <= 16'h0000;
// mem[539] <= 16'h0200;
// mem[540] <= 16'h0200;
// mem[541] <= 16'hf7ff;
// mem[542] <= 16'h0500;
// mem[543] <= 16'h0000;
// mem[544] <= 16'h0000;
// mem[545] <= 16'hfdff;
// mem[546] <= 16'h0200;
// mem[547] <= 16'h0700;
// mem[548] <= 16'h0200;
// mem[549] <= 16'h0000;
// mem[550] <= 16'h0000;
// mem[551] <= 16'h0400;
// mem[552] <= 16'h0200;
// mem[553] <= 16'h0000;
// mem[554] <= 16'h0200;
// mem[555] <= 16'h0300;
// mem[556] <= 16'hfdff;
// mem[557] <= 16'h0900;
// mem[558] <= 16'h0500;
// mem[559] <= 16'h0200;
// mem[560] <= 16'h0400;
// mem[561] <= 16'h0200;
// mem[562] <= 16'h0200;
// mem[563] <= 16'h0200;
// mem[564] <= 16'hfdff;
// mem[565] <= 16'h0200;
// mem[566] <= 16'h0000;
// mem[567] <= 16'hfbff;
// mem[568] <= 16'h0400;
// mem[569] <= 16'h0400;
// mem[570] <= 16'hffff;
// mem[571] <= 16'h0200;
// mem[572] <= 16'h0200;
// mem[573] <= 16'h0200;
// mem[574] <= 16'h0000;
// mem[575] <= 16'h0200;
// mem[576] <= 16'h0200;
// mem[577] <= 16'h0300;
// mem[578] <= 16'h0000;
// mem[579] <= 16'h0300;
// mem[580] <= 16'hfbff;
// mem[581] <= 16'h0200;
// mem[582] <= 16'h0500;
// mem[583] <= 16'h0000;
// mem[584] <= 16'h0300;
// mem[585] <= 16'h0400;
// mem[586] <= 16'hfdff;
// mem[587] <= 16'h0500;
// mem[588] <= 16'hfbff;
// mem[589] <= 16'h0500;
// mem[590] <= 16'h0700;
// mem[591] <= 16'h0200;
// mem[592] <= 16'h0300;
// mem[593] <= 16'hfbff;
// mem[594] <= 16'h0200;
// mem[595] <= 16'h0000;
// mem[596] <= 16'h0000;
// mem[597] <= 16'h0200;
// mem[598] <= 16'h0700;
// mem[599] <= 16'h0000;
// mem[600] <= 16'h0000;
// mem[601] <= 16'h0900;
// mem[602] <= 16'hffff;
// mem[603] <= 16'h0000;
// mem[604] <= 16'h0500;
// mem[605] <= 16'h0200;
// mem[606] <= 16'h0400;
// mem[607] <= 16'h0500;
// mem[608] <= 16'hffff;
// mem[609] <= 16'h0200;
// mem[610] <= 16'h0200;
// mem[611] <= 16'hfbff;
// mem[612] <= 16'h0900;
// mem[613] <= 16'hf9ff;
// mem[614] <= 16'hffff;
// mem[615] <= 16'h0300;
// mem[616] <= 16'hffff;
// mem[617] <= 16'h0400;
// mem[618] <= 16'h0200;
// mem[619] <= 16'h0200;
// mem[620] <= 16'h0300;
// mem[621] <= 16'hffff;
// mem[622] <= 16'h0000;
// mem[623] <= 16'h0500;
// mem[624] <= 16'h0000;
// mem[625] <= 16'h0000;
// mem[626] <= 16'hfdff;
// mem[627] <= 16'hfdff;
// mem[628] <= 16'h0b00;
// mem[629] <= 16'hf9ff;
// mem[630] <= 16'h0300;
// mem[631] <= 16'h0200;
// mem[632] <= 16'h0000;
// mem[633] <= 16'h0200;
// mem[634] <= 16'h0000;
// mem[635] <= 16'h0400;
// mem[636] <= 16'hfdff;
// mem[637] <= 16'h0200;
// mem[638] <= 16'hfbff;
// mem[639] <= 16'hfdff;
// mem[640] <= 16'h0200;
// mem[641] <= 16'hffff;
// mem[642] <= 16'hfdff;
// mem[643] <= 16'h0000;
// mem[644] <= 16'h0000;
// mem[645] <= 16'h0200;
// mem[646] <= 16'hffff;
// mem[647] <= 16'hfdff;
// mem[648] <= 16'hffff;
// mem[649] <= 16'h0200;
// mem[650] <= 16'hf9ff;
// mem[651] <= 16'h0200;
// mem[652] <= 16'h0500;
// mem[653] <= 16'hfbff;
// mem[654] <= 16'h0200;
// mem[655] <= 16'h0000;
// mem[656] <= 16'hffff;
// mem[657] <= 16'hfbff;
// mem[658] <= 16'hfbff;
// mem[659] <= 16'h0300;
// mem[660] <= 16'hf9ff;
// mem[661] <= 16'hf7ff;
// mem[662] <= 16'h0700;
// mem[663] <= 16'hfbff;
// mem[664] <= 16'h0000;
// mem[665] <= 16'hfdff;
// mem[666] <= 16'h0400;
// mem[667] <= 16'hffff;
// mem[668] <= 16'h0000;
// mem[669] <= 16'hf7ff;
// mem[670] <= 16'h0000;
// mem[671] <= 16'h0000;
// mem[672] <= 16'hffff;
// mem[673] <= 16'hffff;
// mem[674] <= 16'hfdff;
// mem[675] <= 16'hfbff;
// mem[676] <= 16'h0000;
// mem[677] <= 16'hfdff;
// mem[678] <= 16'hffff;
// mem[679] <= 16'hfcff;
// mem[680] <= 16'h0000;
// mem[681] <= 16'hfdff;
// mem[682] <= 16'hfbff;
// mem[683] <= 16'h0200;
// mem[684] <= 16'hf9ff;
// mem[685] <= 16'h0000;
// mem[686] <= 16'hffff;
// mem[687] <= 16'hfdff;
// mem[688] <= 16'hfbff;
// mem[689] <= 16'hf9ff;
// mem[690] <= 16'hfdff;
// mem[691] <= 16'hfdff;
// mem[692] <= 16'hfdff;
// mem[693] <= 16'hffff;
// mem[694] <= 16'hfbff;
// mem[695] <= 16'hfbff;
// mem[696] <= 16'hffff;
// mem[697] <= 16'hfeff;
// mem[698] <= 16'hf7ff;
// mem[699] <= 16'hffff;
// mem[700] <= 16'h0300;
// mem[701] <= 16'hfbff;
// mem[702] <= 16'hfdff;
// mem[703] <= 16'hfdff;
// mem[704] <= 16'hfdff;
// mem[705] <= 16'hfdff;
// mem[706] <= 16'hffff;
// mem[707] <= 16'h0000;
// mem[708] <= 16'hfbff;
// mem[709] <= 16'hf3ff;
// mem[710] <= 16'hfdff;
// mem[711] <= 16'hffff;
// mem[712] <= 16'hf7ff;
// mem[713] <= 16'hffff;
// mem[714] <= 16'hfbff;
// mem[715] <= 16'hfdff;
// mem[716] <= 16'h0000;
// mem[717] <= 16'hf5ff;
// mem[718] <= 16'hfeff;
// mem[719] <= 16'h0200;
// mem[720] <= 16'hf7ff;
// mem[721] <= 16'hfdff;
// mem[722] <= 16'hf9ff;
// mem[723] <= 16'hfdff;
// mem[724] <= 16'hfdff;
// mem[725] <= 16'hfbff;
// mem[726] <= 16'hffff;
// mem[727] <= 16'hf5ff;
// mem[728] <= 16'h0400;
// mem[729] <= 16'hffff;
// mem[730] <= 16'hfdff;
// mem[731] <= 16'hfbff;
// mem[732] <= 16'hffff;
// mem[733] <= 16'hffff;
// mem[734] <= 16'hfbff;
// mem[735] <= 16'hf3ff;
// mem[736] <= 16'h0400;
// mem[737] <= 16'hf3ff;
// mem[738] <= 16'hffff;
// mem[739] <= 16'hfdff;
// mem[740] <= 16'hf9ff;
// mem[741] <= 16'hfbff;
// mem[742] <= 16'hfbff;
// mem[743] <= 16'hf7ff;
// mem[744] <= 16'hfbff;
// mem[745] <= 16'hf9ff;
// mem[746] <= 16'hfbff;
// mem[747] <= 16'hfbff;
// mem[748] <= 16'hffff;
// mem[749] <= 16'h0200;
// mem[750] <= 16'hfbff;
// mem[751] <= 16'hffff;
// mem[752] <= 16'hf7ff;
// mem[753] <= 16'hfeff;
// mem[754] <= 16'hffff;
// mem[755] <= 16'hfbff;
// mem[756] <= 16'h0000;
// mem[757] <= 16'hfdff;
// mem[758] <= 16'hfdff;
// mem[759] <= 16'h0200;
// mem[760] <= 16'hf9ff;
// mem[761] <= 16'hf2ff;
// mem[762] <= 16'h0300;
// mem[763] <= 16'hf9ff;
// mem[764] <= 16'hfbff;
// mem[765] <= 16'hfdff;
// mem[766] <= 16'hffff;
// mem[767] <= 16'hfdff;
// mem[768] <= 16'hf9ff;
// mem[769] <= 16'hfbff;
// mem[770] <= 16'hfbff;
// mem[771] <= 16'hffff;
// mem[772] <= 16'hf0ff;
// mem[773] <= 16'hfdff;
// mem[774] <= 16'hfbff;
// mem[775] <= 16'hfbff;
// mem[776] <= 16'hf7ff;
// mem[777] <= 16'hf9ff;
// mem[778] <= 16'hf3ff;
// mem[779] <= 16'hfbff;
// mem[780] <= 16'h0000;
// mem[781] <= 16'hfbff;
// mem[782] <= 16'hffff;
// mem[783] <= 16'hf9ff;
// mem[784] <= 16'hf9ff;
// mem[785] <= 16'hfdff;
// mem[786] <= 16'hfdff;
// mem[787] <= 16'hfbff;
// mem[788] <= 16'hfbff;
// mem[789] <= 16'hf9ff;
// mem[790] <= 16'hfbff;
// mem[791] <= 16'hfdff;
// mem[792] <= 16'hfdff;
// mem[793] <= 16'hf9ff;
// mem[794] <= 16'hfdff;
// mem[795] <= 16'hf5ff;
// mem[796] <= 16'hf2ff;
// mem[797] <= 16'h0000;
// mem[798] <= 16'hfbff;
// mem[799] <= 16'hf9ff;
// mem[800] <= 16'hfdff;
// mem[801] <= 16'hfdff;
// mem[802] <= 16'hf2ff;
// mem[803] <= 16'h0200;
// mem[804] <= 16'hf9ff;
// mem[805] <= 16'hffff;
// mem[806] <= 16'hfbff;
// mem[807] <= 16'hffff;
// mem[808] <= 16'hfdff;
// mem[809] <= 16'hfbff;
// mem[810] <= 16'hfbff;
// mem[811] <= 16'h0000;
// mem[812] <= 16'hf9ff;
// mem[813] <= 16'hf7ff;
// mem[814] <= 16'hf7ff;
// mem[815] <= 16'hf2ff;
// mem[816] <= 16'h0300;
// mem[817] <= 16'hf9ff;
// mem[818] <= 16'hfdff;
// mem[819] <= 16'hf3ff;
// mem[820] <= 16'hf9ff;
// mem[821] <= 16'hfbff;
// mem[822] <= 16'hf7ff;
// mem[823] <= 16'hffff;
// mem[824] <= 16'hfbff;
// mem[825] <= 16'hf7ff;
// mem[826] <= 16'h0000;
// mem[827] <= 16'hfbff;
// mem[828] <= 16'hf9ff;
// mem[829] <= 16'hfbff;
// mem[830] <= 16'hf3ff;
// mem[831] <= 16'h0000;
// mem[832] <= 16'hf7ff;
// mem[833] <= 16'h0200;
// mem[834] <= 16'hffff;
// mem[835] <= 16'hfdff;
// mem[836] <= 16'hfbff;
// mem[837] <= 16'hfbff;
// mem[838] <= 16'hffff;
// mem[839] <= 16'hf9ff;
// mem[840] <= 16'hffff;
// mem[841] <= 16'hfbff;
// mem[842] <= 16'hf9ff;
// mem[843] <= 16'hfbff;
// mem[844] <= 16'hfbff;
// mem[845] <= 16'hfdff;
// mem[846] <= 16'hf9ff;
// mem[847] <= 16'hfdff;
// mem[848] <= 16'hf3ff;
// mem[849] <= 16'h0200;
// mem[850] <= 16'hfbff;
// mem[851] <= 16'hf9ff;
// mem[852] <= 16'hfbff;
// mem[853] <= 16'hfdff;
// mem[854] <= 16'hfbff;
// mem[855] <= 16'hfbff;
// mem[856] <= 16'hfbff;
// mem[857] <= 16'hf7ff;
// mem[858] <= 16'h0200;
// mem[859] <= 16'hf7ff;
// mem[860] <= 16'hfdff;
// mem[861] <= 16'hf4ff;
// mem[862] <= 16'hffff;
// mem[863] <= 16'hffff;
// mem[864] <= 16'hfdff;
// mem[865] <= 16'hffff;
// mem[866] <= 16'hfbff;
// mem[867] <= 16'hffff;
// mem[868] <= 16'hfbff;
// mem[869] <= 16'h0000;
// mem[870] <= 16'hfdff;
// mem[871] <= 16'hfdff;
// mem[872] <= 16'hfdff;
// mem[873] <= 16'hffff;
// mem[874] <= 16'hf4ff;
// mem[875] <= 16'h0200;
// mem[876] <= 16'h0000;
// mem[877] <= 16'hf9ff;
// mem[878] <= 16'hffff;
// mem[879] <= 16'h0000;
// mem[880] <= 16'hfdff;
// mem[881] <= 16'hfbff;
// mem[882] <= 16'h0700;
// mem[883] <= 16'hffff;
// mem[884] <= 16'hffff;
// mem[885] <= 16'h0000;
// mem[886] <= 16'h0000;
// mem[887] <= 16'hffff;
// mem[888] <= 16'hffff;
// mem[889] <= 16'hf5ff;
// mem[890] <= 16'h0400;
// mem[891] <= 16'hffff;
// mem[892] <= 16'hfbff;
// mem[893] <= 16'hffff;
// mem[894] <= 16'h0200;
// mem[895] <= 16'hf5ff;
// mem[896] <= 16'hfdff;
// mem[897] <= 16'h0200;
// mem[898] <= 16'h0000;
// mem[899] <= 16'h0000;
// mem[900] <= 16'h0000;
// mem[901] <= 16'hf9ff;
// mem[902] <= 16'h0000;
// mem[903] <= 16'h0500;
// mem[904] <= 16'hf7ff;
// mem[905] <= 16'h0200;
// mem[906] <= 16'hf7ff;
// mem[907] <= 16'hffff;
// mem[908] <= 16'h0300;
// mem[909] <= 16'hffff;
// mem[910] <= 16'hfdff;
// mem[911] <= 16'h0200;
// mem[912] <= 16'h0200;
// mem[913] <= 16'h0300;
// mem[914] <= 16'h0500;
// mem[915] <= 16'hffff;
// mem[916] <= 16'h0500;
// mem[917] <= 16'h0000;
// mem[918] <= 16'h0200;
// mem[919] <= 16'hffff;
// mem[920] <= 16'h0500;
// mem[921] <= 16'hfbff;
// mem[922] <= 16'h0200;
// mem[923] <= 16'h0300;
// mem[924] <= 16'hffff;
// mem[925] <= 16'h0400;
// mem[926] <= 16'h0000;
// mem[927] <= 16'h0300;
// mem[928] <= 16'h0000;
// mem[929] <= 16'h0400;
// mem[930] <= 16'hf7ff;
// mem[931] <= 16'h0900;
// mem[932] <= 16'h0200;
// mem[933] <= 16'hffff;
// mem[934] <= 16'h0500;
// mem[935] <= 16'h0000;
// mem[936] <= 16'h0200;
// mem[937] <= 16'h0200;
// mem[938] <= 16'h0200;
// mem[939] <= 16'h0700;
// mem[940] <= 16'h0200;
// mem[941] <= 16'h0300;
// mem[942] <= 16'h0300;
// mem[943] <= 16'h0200;
// mem[944] <= 16'hfbff;
// mem[945] <= 16'h0900;
// mem[946] <= 16'h0300;
// mem[947] <= 16'h0400;
// mem[948] <= 16'h0200;
// mem[949] <= 16'h0700;
// mem[950] <= 16'h0300;
// mem[951] <= 16'h0500;
// mem[952] <= 16'h0000;
// mem[953] <= 16'h0500;
// mem[954] <= 16'hfdff;
// mem[955] <= 16'h0200;
// mem[956] <= 16'h0b00;
// mem[957] <= 16'h0200;
// mem[958] <= 16'h0500;
// mem[959] <= 16'h0000;
// mem[960] <= 16'h0500;
// mem[961] <= 16'h0200;
// mem[962] <= 16'h0500;
// mem[963] <= 16'h0500;
// mem[964] <= 16'hffff;
// mem[965] <= 16'h0b00;
// mem[966] <= 16'h0700;
// mem[967] <= 16'h0500;
// mem[968] <= 16'h0700;
// mem[969] <= 16'h0300;
// mem[970] <= 16'h0700;
// mem[971] <= 16'h0500;
// mem[972] <= 16'h0700;
// mem[973] <= 16'h0700;
// mem[974] <= 16'h0700;
// mem[975] <= 16'h0400;
// mem[976] <= 16'h0900;
// mem[977] <= 16'h0000;
// mem[978] <= 16'h0700;
// mem[979] <= 16'h0500;
// mem[980] <= 16'h0900;
// mem[981] <= 16'h0b00;
// mem[982] <= 16'h0300;
// mem[983] <= 16'h0700;
// mem[984] <= 16'h0500;
// mem[985] <= 16'h0200;
// mem[986] <= 16'h0500;
// mem[987] <= 16'h0300;
// mem[988] <= 16'h0000;
// mem[989] <= 16'h0d00;
// mem[990] <= 16'h0500;
// mem[991] <= 16'h0300;
// mem[992] <= 16'h0200;
// mem[993] <= 16'h0500;
// mem[994] <= 16'h0400;
// mem[995] <= 16'h0700;
// mem[996] <= 16'h0300;
// mem[997] <= 16'h0500;
// mem[998] <= 16'h0300;
// mem[999] <= 16'h0500;
// mem[1000] <= 16'h0000;
// mem[1001] <= 16'h0900;
// mem[1002] <= 16'h0000;
// mem[1003] <= 16'h0200;
// mem[1004] <= 16'h0500;
// mem[1005] <= 16'h0200;
// mem[1006] <= 16'h0900;
// mem[1007] <= 16'hfdff;
// mem[1008] <= 16'h0b00;
// mem[1009] <= 16'h0300;
// mem[1010] <= 16'h0500;
// mem[1011] <= 16'h0400;
// mem[1012] <= 16'h0200;
// mem[1013] <= 16'h0300;
// mem[1014] <= 16'hfdff;
// mem[1015] <= 16'h0f00;
// mem[1016] <= 16'hfbff;
// mem[1017] <= 16'h0300;
// mem[1018] <= 16'h0900;
// mem[1019] <= 16'h0300;
// mem[1020] <= 16'h0000;
// mem[1021] <= 16'h0500;
// mem[1022] <= 16'hfdff;
// mem[1023] <= 16'h0b00;
// mem[1024] <= 16'hfbff;
// mem[1025] <= 16'h0700;
// mem[1026] <= 16'h0200;
// mem[1027] <= 16'h0000;
// mem[1028] <= 16'h0b00;
// mem[1029] <= 16'h0000;
// mem[1030] <= 16'h0200;
// mem[1031] <= 16'h0200;
// mem[1032] <= 16'h0200;
// mem[1033] <= 16'hfdff;
// mem[1034] <= 16'hf9ff;
// mem[1035] <= 16'h0f00;
// mem[1036] <= 16'hfbff;
// mem[1037] <= 16'h0200;
// mem[1038] <= 16'h0700;
// mem[1039] <= 16'hffff;
// mem[1040] <= 16'hffff;
// mem[1041] <= 16'h0200;
// mem[1042] <= 16'hfbff;
// mem[1043] <= 16'h0200;
// mem[1044] <= 16'h0200;
// mem[1045] <= 16'hffff;
// mem[1046] <= 16'h0200;
// mem[1047] <= 16'h0000;
// mem[1048] <= 16'h0000;
// mem[1049] <= 16'h0000;
// mem[1050] <= 16'h0200;
// mem[1051] <= 16'hf7ff;
// mem[1052] <= 16'h0300;
// mem[1053] <= 16'h0400;
// mem[1054] <= 16'hffff;
// mem[1055] <= 16'hf9ff;
// mem[1056] <= 16'h0900;
// mem[1057] <= 16'h0500;
// mem[1058] <= 16'h0300;
// mem[1059] <= 16'hffff;
// mem[1060] <= 16'hfeff;
// mem[1061] <= 16'h0000;
// mem[1062] <= 16'hffff;
// mem[1063] <= 16'h0000;
// mem[1064] <= 16'h0000;
// mem[1065] <= 16'h0200;
// mem[1066] <= 16'hf9ff;
// mem[1067] <= 16'h0700;
// mem[1068] <= 16'hffff;
// mem[1069] <= 16'hfdff;
// mem[1070] <= 16'h0900;
// mem[1071] <= 16'hffff;
// mem[1072] <= 16'h0400;
// mem[1073] <= 16'hf9ff;
// mem[1074] <= 16'h0500;
// mem[1075] <= 16'h0200;
// mem[1076] <= 16'hfdff;
// mem[1077] <= 16'h0400;
// mem[1078] <= 16'hf5ff;
// mem[1079] <= 16'h0200;
// mem[1080] <= 16'h0400;
// mem[1081] <= 16'h0000;
// mem[1082] <= 16'hfdff;
// mem[1083] <= 16'h0400;
// mem[1084] <= 16'hfbff;
// mem[1085] <= 16'h0000;
// mem[1086] <= 16'hfbff;
// mem[1087] <= 16'h0000;
// mem[1088] <= 16'hfbff;
// mem[1089] <= 16'hf7ff;
// mem[1090] <= 16'h0500;
// mem[1091] <= 16'h0200;
// mem[1092] <= 16'hf9ff;
// mem[1093] <= 16'hfdff;
// mem[1094] <= 16'h0500;
// mem[1095] <= 16'hf9ff;
// mem[1096] <= 16'h0500;
// mem[1097] <= 16'hf3ff;
// mem[1098] <= 16'hffff;
// mem[1099] <= 16'h0000;
// mem[1100] <= 16'h0000;
// mem[1101] <= 16'hf9ff;
// mem[1102] <= 16'h0600;
// mem[1103] <= 16'hfdff;
// mem[1104] <= 16'hffff;
// mem[1105] <= 16'h0500;
// mem[1106] <= 16'hffff;
// mem[1107] <= 16'h0000;
// mem[1108] <= 16'hffff;
// mem[1109] <= 16'hfbff;
// mem[1110] <= 16'hffff;
// mem[1111] <= 16'hf9ff;
// mem[1112] <= 16'hffff;
// mem[1113] <= 16'h0400;
// mem[1114] <= 16'hf3ff;
// mem[1115] <= 16'h0200;
// mem[1116] <= 16'hfdff;
// mem[1117] <= 16'hfdff;
// mem[1118] <= 16'hfdff;
// mem[1119] <= 16'hffff;
// mem[1120] <= 16'hffff;
// mem[1121] <= 16'hfdff;
// mem[1122] <= 16'hfdff;
// mem[1123] <= 16'hfdff;
// mem[1124] <= 16'hffff;
// mem[1125] <= 16'hf7ff;
// mem[1126] <= 16'hfbff;
// mem[1127] <= 16'hffff;
// mem[1128] <= 16'hffff;
// mem[1129] <= 16'h0000;
// mem[1130] <= 16'hffff;
// mem[1131] <= 16'hf9ff;
// mem[1132] <= 16'h0200;
// mem[1133] <= 16'hf1ff;
// mem[1134] <= 16'hffff;
// mem[1135] <= 16'hfdff;
// mem[1136] <= 16'hf9ff;
// mem[1137] <= 16'h0200;
// mem[1138] <= 16'hfdff;
// mem[1139] <= 16'hfdff;
// mem[1140] <= 16'hfdff;
// mem[1141] <= 16'h0300;
// mem[1142] <= 16'heeff;
// mem[1143] <= 16'h0300;
// mem[1144] <= 16'hf5ff;
// mem[1145] <= 16'hfbff;
// mem[1146] <= 16'h0300;
// mem[1147] <= 16'hf1ff;
// mem[1148] <= 16'h0000;
// mem[1149] <= 16'hf7ff;
// mem[1150] <= 16'h0700;
// mem[1151] <= 16'hf9ff;
// mem[1152] <= 16'hf9ff;
// mem[1153] <= 16'hfbff;
// mem[1154] <= 16'hfbff;
// mem[1155] <= 16'h0000;
// mem[1156] <= 16'hf0ff;
// mem[1157] <= 16'h0700;
// mem[1158] <= 16'hf2ff;
// mem[1159] <= 16'hffff;
// mem[1160] <= 16'hf9ff;
// mem[1161] <= 16'h0000;
// mem[1162] <= 16'h0300;
// mem[1163] <= 16'hf3ff;
// mem[1164] <= 16'h0400;
// mem[1165] <= 16'hf7ff;
// mem[1166] <= 16'hffff;
// mem[1167] <= 16'h0400;
// mem[1168] <= 16'hf2ff;
// mem[1169] <= 16'h0200;
// mem[1170] <= 16'hf9ff;
// mem[1171] <= 16'hf9ff;
// mem[1172] <= 16'h0200;
// mem[1173] <= 16'hfbff;
// mem[1174] <= 16'hffff;
// mem[1175] <= 16'hfbff;
// mem[1176] <= 16'hfdff;
// mem[1177] <= 16'hf1ff;
// mem[1178] <= 16'h0500;
// mem[1179] <= 16'hf9ff;
// mem[1180] <= 16'h0000;
// mem[1181] <= 16'hf5ff;
// mem[1182] <= 16'hfdff;
// mem[1183] <= 16'hffff;
// mem[1184] <= 16'hfdff;
// mem[1185] <= 16'hf9ff;
// mem[1186] <= 16'hfdff;
// mem[1187] <= 16'hf5ff;
// mem[1188] <= 16'hffff;
// mem[1189] <= 16'hffff;
// mem[1190] <= 16'hf3ff;
// mem[1191] <= 16'h0400;
// mem[1192] <= 16'hfdff;
// mem[1193] <= 16'hfbff;
// mem[1194] <= 16'hfdff;
// mem[1195] <= 16'hf7ff;
// mem[1196] <= 16'h0000;
// mem[1197] <= 16'hffff;
// mem[1198] <= 16'hf5ff;
// mem[1199] <= 16'hfbff;
// mem[1200] <= 16'h0000;
// mem[1201] <= 16'hf9ff;
// mem[1202] <= 16'hfbff;
// mem[1203] <= 16'hfeff;
// mem[1204] <= 16'hfdff;
// mem[1205] <= 16'hfbff;
// mem[1206] <= 16'hffff;
// mem[1207] <= 16'hffff;
// mem[1208] <= 16'hfbff;
// mem[1209] <= 16'hfbff;
// mem[1210] <= 16'hfbff;
// mem[1211] <= 16'hf3ff;
// mem[1212] <= 16'hffff;
// mem[1213] <= 16'hf7ff;
// mem[1214] <= 16'hfbff;
// mem[1215] <= 16'hfdff;
// mem[1216] <= 16'hfbff;
// mem[1217] <= 16'hf7ff;
// mem[1218] <= 16'hffff;
// mem[1219] <= 16'hf7ff;
// mem[1220] <= 16'hfbff;
// mem[1221] <= 16'hf9ff;
// mem[1222] <= 16'hfdff;
// mem[1223] <= 16'hfbff;
// mem[1224] <= 16'hf5ff;
// mem[1225] <= 16'hfdff;
// mem[1226] <= 16'hfdff;
// mem[1227] <= 16'hfbff;
// mem[1228] <= 16'hf9ff;
// mem[1229] <= 16'hf9ff;
// mem[1230] <= 16'hf9ff;
// mem[1231] <= 16'hf9ff;
// mem[1232] <= 16'hfbff;
// mem[1233] <= 16'hf7ff;
// mem[1234] <= 16'hf7ff;
// mem[1235] <= 16'h0000;
// mem[1236] <= 16'hf5ff;
// mem[1237] <= 16'hfbff;
// mem[1238] <= 16'hf3ff;
// mem[1239] <= 16'hfdff;
// mem[1240] <= 16'hf2ff;
// mem[1241] <= 16'hf9ff;
// mem[1242] <= 16'hfbff;
// mem[1243] <= 16'hf9ff;
// mem[1244] <= 16'hfbff;
// mem[1245] <= 16'hf9ff;
// mem[1246] <= 16'hf9ff;
// mem[1247] <= 16'hfbff;
// mem[1248] <= 16'hffff;
// mem[1249] <= 16'hf7ff;
// mem[1250] <= 16'hfbff;
// mem[1251] <= 16'hf7ff;
// mem[1252] <= 16'hf7ff;
// mem[1253] <= 16'hfbff;
// mem[1254] <= 16'hf5ff;
// mem[1255] <= 16'h0500;
// mem[1256] <= 16'hecff;
// mem[1257] <= 16'h0200;
// mem[1258] <= 16'hffff;
// mem[1259] <= 16'hf0ff;
// mem[1260] <= 16'h0900;
// mem[1261] <= 16'heeff;
// mem[1262] <= 16'hfdff;
// mem[1263] <= 16'hf7ff;
// mem[1264] <= 16'h0000;
// mem[1265] <= 16'hf7ff;
// mem[1266] <= 16'hf9ff;
// mem[1267] <= 16'hfbff;
// mem[1268] <= 16'hf9ff;
// mem[1269] <= 16'hf9ff;
// mem[1270] <= 16'hfdff;
// mem[1271] <= 16'hf5ff;
// mem[1272] <= 16'h0000;
// mem[1273] <= 16'hf9ff;
// mem[1274] <= 16'hfbff;
// mem[1275] <= 16'hfeff;
// mem[1276] <= 16'hf3ff;
// mem[1277] <= 16'h0200;
// mem[1278] <= 16'heeff;
// mem[1279] <= 16'h0300;
// mem[1280] <= 16'hf3ff;
// mem[1281] <= 16'hfbff;
// mem[1282] <= 16'hf7ff;
// mem[1283] <= 16'hf9ff;
// mem[1284] <= 16'hf9ff;
// mem[1285] <= 16'hf0ff;
// mem[1286] <= 16'h0200;
// mem[1287] <= 16'hf9ff;
// mem[1288] <= 16'h0200;
// mem[1289] <= 16'hf0ff;
// mem[1290] <= 16'hffff;
// mem[1291] <= 16'h0200;
// mem[1292] <= 16'hf7ff;
// mem[1293] <= 16'hfbff;
// mem[1294] <= 16'hf9ff;
// mem[1295] <= 16'hf9ff;
// mem[1296] <= 16'h0500;
// mem[1297] <= 16'hf7ff;
// mem[1298] <= 16'hfdff;
// mem[1299] <= 16'hf7ff;
// mem[1300] <= 16'h0300;
// mem[1301] <= 16'hfdff;
// mem[1302] <= 16'hfbff;
// mem[1303] <= 16'h0200;
// mem[1304] <= 16'hf7ff;
// mem[1305] <= 16'hffff;
// mem[1306] <= 16'hfdff;
// mem[1307] <= 16'hfbff;
// mem[1308] <= 16'h0000;
// mem[1309] <= 16'hf9ff;
// mem[1310] <= 16'h0000;
// mem[1311] <= 16'hfbff;
// mem[1312] <= 16'hfdff;
// mem[1313] <= 16'hf9ff;
// mem[1314] <= 16'hf9ff;
// mem[1315] <= 16'h0200;
// mem[1316] <= 16'hfbff;
// mem[1317] <= 16'hf9ff;
// mem[1318] <= 16'hfbff;
// mem[1319] <= 16'h0500;
// mem[1320] <= 16'hfbff;
// mem[1321] <= 16'h0200;
// mem[1322] <= 16'hf5ff;
// mem[1323] <= 16'h0200;
// mem[1324] <= 16'h0700;
// mem[1325] <= 16'hffff;
// mem[1326] <= 16'h0200;
// mem[1327] <= 16'hffff;
// mem[1328] <= 16'h0500;
// mem[1329] <= 16'hfdff;
// mem[1330] <= 16'h0000;
// mem[1331] <= 16'h0400;
// mem[1332] <= 16'hffff;
// mem[1333] <= 16'h0600;
// mem[1334] <= 16'h0000;
// mem[1335] <= 16'h0300;
// mem[1336] <= 16'hfdff;
// mem[1337] <= 16'h0000;
// mem[1338] <= 16'h0700;
// mem[1339] <= 16'h0000;
// mem[1340] <= 16'h0300;
// mem[1341] <= 16'hffff;
// mem[1342] <= 16'hfdff;
// mem[1343] <= 16'h0000;
// mem[1344] <= 16'h0200;
// mem[1345] <= 16'hffff;
// mem[1346] <= 16'h0200;
// mem[1347] <= 16'h0000;
// mem[1348] <= 16'h0300;
// mem[1349] <= 16'h0400;
// mem[1350] <= 16'h0400;
// mem[1351] <= 16'h0300;
// mem[1352] <= 16'h0200;
// mem[1353] <= 16'h0200;
// mem[1354] <= 16'h0300;
// mem[1355] <= 16'h0700;
// mem[1356] <= 16'h0300;
// mem[1357] <= 16'h0700;
// mem[1358] <= 16'hfbff;
// mem[1359] <= 16'h0700;
// mem[1360] <= 16'h0700;
// mem[1361] <= 16'h0200;
// mem[1362] <= 16'h0700;
// mem[1363] <= 16'hfdff;
// mem[1364] <= 16'h0200;
// mem[1365] <= 16'h0300;
// mem[1366] <= 16'h0000;
// mem[1367] <= 16'h0500;
// mem[1368] <= 16'h0300;
// mem[1369] <= 16'h0200;
// mem[1370] <= 16'h0000;
// mem[1371] <= 16'h0200;
// mem[1372] <= 16'h0000;
// mem[1373] <= 16'h0500;
// mem[1374] <= 16'h0200;
// mem[1375] <= 16'hf9ff;
// mem[1376] <= 16'h0300;
// mem[1377] <= 16'h0000;
// mem[1378] <= 16'h0700;
// mem[1379] <= 16'h0300;
// mem[1380] <= 16'h0900;
// mem[1381] <= 16'h0200;
// mem[1382] <= 16'h0500;
// mem[1383] <= 16'hfdff;
// mem[1384] <= 16'h0000;
// mem[1385] <= 16'h0b00;
// mem[1386] <= 16'h0300;
// mem[1387] <= 16'h0500;
// mem[1388] <= 16'hf7ff;
// mem[1389] <= 16'h0f00;
// mem[1390] <= 16'hffff;
// mem[1391] <= 16'h0200;
// mem[1392] <= 16'h0700;
// mem[1393] <= 16'hf7ff;
// mem[1394] <= 16'h0700;
// mem[1395] <= 16'hffff;
// mem[1396] <= 16'h0900;
// mem[1397] <= 16'hffff;
// mem[1398] <= 16'hffff;
// mem[1399] <= 16'h0d00;
// mem[1400] <= 16'hfbff;
// mem[1401] <= 16'h0d00;
// mem[1402] <= 16'hffff;
// mem[1403] <= 16'hfdff;
// mem[1404] <= 16'h0400;
// mem[1405] <= 16'h0000;
// mem[1406] <= 16'h0900;
// mem[1407] <= 16'hf3ff;
// mem[1408] <= 16'h0f00;
// mem[1409] <= 16'hffff;
// mem[1410] <= 16'h0000;
// mem[1411] <= 16'h0300;
// mem[1412] <= 16'hfdff;
// mem[1413] <= 16'h0500;
// mem[1414] <= 16'hf7ff;
// mem[1415] <= 16'h0f00;
// mem[1416] <= 16'hfbff;
// mem[1417] <= 16'h0200;
// mem[1418] <= 16'h0300;
// mem[1419] <= 16'h0200;
// mem[1420] <= 16'h0200;
// mem[1421] <= 16'hf9ff;
// mem[1422] <= 16'h0000;
// mem[1423] <= 16'hfeff;
// mem[1424] <= 16'hffff;
// mem[1425] <= 16'hfbff;
// mem[1426] <= 16'hfdff;
// mem[1427] <= 16'h0300;
// mem[1428] <= 16'h0500;
// mem[1429] <= 16'hf7ff;
// mem[1430] <= 16'h0700;
// mem[1431] <= 16'hf9ff;
// mem[1432] <= 16'h0000;
// mem[1433] <= 16'h0700;
// mem[1434] <= 16'h0000;
// mem[1435] <= 16'hfdff;
// mem[1436] <= 16'hf7ff;
// mem[1437] <= 16'h0400;
// mem[1438] <= 16'hfdff;
// mem[1439] <= 16'hfdff;
// mem[1440] <= 16'h0300;
// mem[1441] <= 16'h0400;
// mem[1442] <= 16'h0000;
// mem[1443] <= 16'hfdff;
// mem[1444] <= 16'h0000;
// mem[1445] <= 16'hfdff;
// mem[1446] <= 16'h0000;
// mem[1447] <= 16'h0300;
// mem[1448] <= 16'h0000;
// mem[1449] <= 16'h0200;
// mem[1450] <= 16'hfdff;
// mem[1451] <= 16'h0500;
// mem[1452] <= 16'h0300;
// mem[1453] <= 16'hfbff;
// mem[1454] <= 16'h0000;
// mem[1455] <= 16'h0500;
// mem[1456] <= 16'hfdff;
// mem[1457] <= 16'hfbff;
// mem[1458] <= 16'h0400;
// mem[1459] <= 16'h0000;
// mem[1460] <= 16'h0000;
// mem[1461] <= 16'hffff;
// mem[1462] <= 16'hfdff;
// mem[1463] <= 16'h0900;
// mem[1464] <= 16'hfbff;
// mem[1465] <= 16'hfdff;
// mem[1466] <= 16'h0000;
// mem[1467] <= 16'hfdff;
// mem[1468] <= 16'h0300;
// mem[1469] <= 16'hf5ff;
// mem[1470] <= 16'h0600;
// mem[1471] <= 16'hfdff;
// mem[1472] <= 16'h0000;
// mem[1473] <= 16'hf9ff;
// mem[1474] <= 16'hfdff;
// mem[1475] <= 16'hfbff;
// mem[1476] <= 16'hfbff;
// mem[1477] <= 16'h0000;
// mem[1478] <= 16'h0000;
// mem[1479] <= 16'h0000;
// mem[1480] <= 16'h0000;
// mem[1481] <= 16'hffff;
// mem[1482] <= 16'h0000;
// mem[1483] <= 16'hfdff;
// mem[1484] <= 16'hfbff;
// mem[1485] <= 16'h0500;
// mem[1486] <= 16'hf9ff;
// mem[1487] <= 16'h0000;
// mem[1488] <= 16'hffff;
// mem[1489] <= 16'h0000;
// mem[1490] <= 16'hf5ff;
// mem[1491] <= 16'h0200;
// mem[1492] <= 16'hfdff;
// mem[1493] <= 16'hfdff;
// mem[1494] <= 16'hfdff;
// mem[1495] <= 16'h0000;
// mem[1496] <= 16'h0200;
// mem[1497] <= 16'h0000;
// mem[1498] <= 16'hffff;
// mem[1499] <= 16'h0000;
// mem[1500] <= 16'hf1ff;
// mem[1501] <= 16'h0200;
// mem[1502] <= 16'h0200;
// mem[1503] <= 16'hf5ff;
// mem[1504] <= 16'h0200;
// mem[1505] <= 16'h0200;
// mem[1506] <= 16'hffff;
// mem[1507] <= 16'h0000;
// mem[1508] <= 16'hf7ff;
// mem[1509] <= 16'h0500;
// mem[1510] <= 16'h0200;
// mem[1511] <= 16'hf7ff;
// mem[1512] <= 16'h0200;
// mem[1513] <= 16'hfdff;
// mem[1514] <= 16'hffff;
// mem[1515] <= 16'h0300;
// mem[1516] <= 16'hffff;
// mem[1517] <= 16'h0200;
// mem[1518] <= 16'hfbff;
// mem[1519] <= 16'h0200;
// mem[1520] <= 16'hfbff;
// mem[1521] <= 16'h0200;
// mem[1522] <= 16'h0200;
// mem[1523] <= 16'hfbff;
// mem[1524] <= 16'hfdff;
// mem[1525] <= 16'h0200;
// mem[1526] <= 16'hfdff;
// mem[1527] <= 16'hf9ff;
// mem[1528] <= 16'h0500;
// mem[1529] <= 16'hf3ff;
// mem[1530] <= 16'h0200;
// mem[1531] <= 16'hfbff;
// mem[1532] <= 16'hfdff;
// mem[1533] <= 16'hf7ff;
// mem[1534] <= 16'hfbff;
// mem[1535] <= 16'hfdff;
// mem[1536] <= 16'hf9ff;
// mem[1537] <= 16'hf0ff;
// mem[1538] <= 16'h0200;
// mem[1539] <= 16'h0000;
// mem[1540] <= 16'hffff;
// mem[1541] <= 16'hffff;
// mem[1542] <= 16'hffff;
// mem[1543] <= 16'h0200;
// mem[1544] <= 16'hf5ff;
// mem[1545] <= 16'h0200;
// mem[1546] <= 16'hfdff;
// mem[1547] <= 16'hfbff;
// mem[1548] <= 16'h0000;
// mem[1549] <= 16'hf5ff;
// mem[1550] <= 16'h0200;
// mem[1551] <= 16'h0200;
// mem[1552] <= 16'hfbff;
// mem[1553] <= 16'hfeff;
// mem[1554] <= 16'hffff;
// mem[1555] <= 16'hfbff;
// mem[1556] <= 16'hfbff;
// mem[1557] <= 16'hffff;
// mem[1558] <= 16'hfbff;
// mem[1559] <= 16'hf9ff;
// mem[1560] <= 16'hffff;
// mem[1561] <= 16'h0000;
// mem[1562] <= 16'hfbff;
// mem[1563] <= 16'hffff;
// mem[1564] <= 16'hf1ff;
// mem[1565] <= 16'h0200;
// mem[1566] <= 16'hfdff;
// mem[1567] <= 16'hf9ff;
// mem[1568] <= 16'hfdff;
// mem[1569] <= 16'hffff;
// mem[1570] <= 16'hfbff;
// mem[1571] <= 16'hfdff;
// mem[1572] <= 16'hfdff;
// mem[1573] <= 16'hffff;
// mem[1574] <= 16'hf7ff;
// mem[1575] <= 16'hf9ff;
// mem[1576] <= 16'h0300;
// mem[1577] <= 16'hfbff;
// mem[1578] <= 16'hfbff;
// mem[1579] <= 16'hf9ff;
// mem[1580] <= 16'hfdff;
// mem[1581] <= 16'hf7ff;
// mem[1582] <= 16'hfbff;
// mem[1583] <= 16'hfbff;
// mem[1584] <= 16'hfeff;
// mem[1585] <= 16'hf7ff;
// mem[1586] <= 16'hf7ff;
// mem[1587] <= 16'h0400;
// mem[1588] <= 16'hfbff;
// mem[1589] <= 16'hf9ff;
// mem[1590] <= 16'hfbff;
// mem[1591] <= 16'hfdff;
// mem[1592] <= 16'hfbff;
// mem[1593] <= 16'hfbff;
// mem[1594] <= 16'hf9ff;
// mem[1595] <= 16'hf7ff;
// mem[1596] <= 16'h0000;
// mem[1597] <= 16'hf5ff;
// mem[1598] <= 16'hfeff;
// mem[1599] <= 16'hf7ff;
// mem[1600] <= 16'hf1ff;
// mem[1601] <= 16'h0000;
// mem[1602] <= 16'hf9ff;
// mem[1603] <= 16'hf9ff;
// mem[1604] <= 16'hfdff;
// mem[1605] <= 16'hfbff;
// mem[1606] <= 16'h0000;
// mem[1607] <= 16'hffff;
// mem[1608] <= 16'hfdff;
// mem[1609] <= 16'hfdff;
// mem[1610] <= 16'hffff;
// mem[1611] <= 16'hf0ff;
// mem[1612] <= 16'h0000;
// mem[1613] <= 16'hfdff;
// mem[1614] <= 16'hf3ff;
// mem[1615] <= 16'h0800;
// mem[1616] <= 16'hf0ff;
// mem[1617] <= 16'h0000;
// mem[1618] <= 16'hfbff;
// mem[1619] <= 16'hffff;
// mem[1620] <= 16'hf7ff;
// mem[1621] <= 16'hf3ff;
// mem[1622] <= 16'h0200;
// mem[1623] <= 16'hf7ff;
// mem[1624] <= 16'hfdff;
// mem[1625] <= 16'hf9ff;
// mem[1626] <= 16'heeff;
// mem[1627] <= 16'h0000;
// mem[1628] <= 16'hf5ff;
// mem[1629] <= 16'hfdff;
// mem[1630] <= 16'hf7ff;
// mem[1631] <= 16'hfbff;
// mem[1632] <= 16'hfdff;
// mem[1633] <= 16'heeff;
// mem[1634] <= 16'h0700;
// mem[1635] <= 16'hf2ff;
// mem[1636] <= 16'hfdff;
// mem[1637] <= 16'hf9ff;
// mem[1638] <= 16'hfdff;
// mem[1639] <= 16'hfbff;
// mem[1640] <= 16'hfdff;
// mem[1641] <= 16'hf9ff;
// mem[1642] <= 16'hfbff;
// mem[1643] <= 16'hffff;
// mem[1644] <= 16'hf7ff;
// mem[1645] <= 16'hfdff;
// mem[1646] <= 16'h0200;
// mem[1647] <= 16'hf5ff;
// mem[1648] <= 16'h0300;
// mem[1649] <= 16'hf3ff;
// mem[1650] <= 16'hf9ff;
// mem[1651] <= 16'h0300;
// mem[1652] <= 16'hf9ff;
// mem[1653] <= 16'hffff;
// mem[1654] <= 16'hf9ff;
// mem[1655] <= 16'hfbff;
// mem[1656] <= 16'hfdff;
// mem[1657] <= 16'hffff;
// mem[1658] <= 16'h0400;
// mem[1659] <= 16'hf3ff;
// mem[1660] <= 16'hffff;
// mem[1661] <= 16'hf9ff;
// mem[1662] <= 16'h0000;
// mem[1663] <= 16'hf7ff;
// mem[1664] <= 16'h0300;
// mem[1665] <= 16'hf0ff;
// mem[1666] <= 16'h0200;
// mem[1667] <= 16'hfdff;
// mem[1668] <= 16'hf7ff;
// mem[1669] <= 16'h0500;
// mem[1670] <= 16'hf3ff;
// mem[1671] <= 16'hf9ff;
// mem[1672] <= 16'h0400;
// mem[1673] <= 16'hf5ff;
// mem[1674] <= 16'h0500;
// mem[1675] <= 16'hf7ff;
// mem[1676] <= 16'h0200;
// mem[1677] <= 16'hf7ff;
// mem[1678] <= 16'hffff;
// mem[1679] <= 16'hffff;
// mem[1680] <= 16'hf9ff;
// mem[1681] <= 16'hfdff;
// mem[1682] <= 16'hf5ff;
// mem[1683] <= 16'h0200;
// mem[1684] <= 16'hfdff;
// mem[1685] <= 16'hfdff;
// mem[1686] <= 16'hfbff;
// mem[1687] <= 16'hf5ff;
// mem[1688] <= 16'h0500;
// mem[1689] <= 16'hf5ff;
// mem[1690] <= 16'hfdff;
// mem[1691] <= 16'h0200;
// mem[1692] <= 16'hfbff;
// mem[1693] <= 16'h0400;
// mem[1694] <= 16'hf5ff;
// mem[1695] <= 16'h0700;
// mem[1696] <= 16'hfdff;
// mem[1697] <= 16'h0200;
// mem[1698] <= 16'h0000;
// mem[1699] <= 16'hfbff;
// mem[1700] <= 16'h0000;
// mem[1701] <= 16'h0000;
// mem[1702] <= 16'hf9ff;
// mem[1703] <= 16'hf9ff;
// mem[1704] <= 16'hffff;
// mem[1705] <= 16'hf9ff;
// mem[1706] <= 16'h0000;
// mem[1707] <= 16'hffff;
// mem[1708] <= 16'h0200;
// mem[1709] <= 16'hffff;
// mem[1710] <= 16'h0000;
// mem[1711] <= 16'hfdff;
// mem[1712] <= 16'h0200;
// mem[1713] <= 16'hffff;
// mem[1714] <= 16'h0200;
// mem[1715] <= 16'hffff;
// mem[1716] <= 16'h0000;
// mem[1717] <= 16'h0200;
// mem[1718] <= 16'h0000;
// mem[1719] <= 16'h0000;
// mem[1720] <= 16'hffff;
// mem[1721] <= 16'hfdff;
// mem[1722] <= 16'h0300;
// mem[1723] <= 16'h0400;
// mem[1724] <= 16'hffff;
// mem[1725] <= 16'h0200;
// mem[1726] <= 16'hf7ff;
// mem[1727] <= 16'h0000;
// mem[1728] <= 16'h0700;
// mem[1729] <= 16'h0000;
// mem[1730] <= 16'hfdff;
// mem[1731] <= 16'h0000;
// mem[1732] <= 16'h0000;
// mem[1733] <= 16'h0300;
// mem[1734] <= 16'h0200;
// mem[1735] <= 16'hfbff;
// mem[1736] <= 16'h0900;
// mem[1737] <= 16'h0000;
// mem[1738] <= 16'h0000;
// mem[1739] <= 16'h0200;
// mem[1740] <= 16'hfbff;
// mem[1741] <= 16'h0200;
// mem[1742] <= 16'h0500;
// mem[1743] <= 16'h0200;
// mem[1744] <= 16'h0300;
// mem[1745] <= 16'h0200;
// mem[1746] <= 16'h0500;
// mem[1747] <= 16'hfbff;
// mem[1748] <= 16'h0900;
// mem[1749] <= 16'h0400;
// mem[1750] <= 16'h0000;
// mem[1751] <= 16'h0900;
// mem[1752] <= 16'h0200;
// mem[1753] <= 16'h0400;
// mem[1754] <= 16'h0300;
// mem[1755] <= 16'h0500;
// mem[1756] <= 16'hfdff;
// mem[1757] <= 16'h0900;
// mem[1758] <= 16'h0200;
// mem[1759] <= 16'h0200;
// mem[1760] <= 16'h0200;
// mem[1761] <= 16'h0500;
// mem[1762] <= 16'h0700;
// mem[1763] <= 16'hfdff;
// mem[1764] <= 16'h0900;
// mem[1765] <= 16'h0300;
// mem[1766] <= 16'h0700;
// mem[1767] <= 16'h0400;
// mem[1768] <= 16'h0300;
// mem[1769] <= 16'h0400;
// mem[1770] <= 16'hffff;
// mem[1771] <= 16'h0d00;
// mem[1772] <= 16'h0700;
// mem[1773] <= 16'h0900;
// mem[1774] <= 16'h0700;
// mem[1775] <= 16'h0500;
// mem[1776] <= 16'h0000;
// mem[1777] <= 16'h0d00;
// mem[1778] <= 16'h0900;
// mem[1779] <= 16'h0000;
// mem[1780] <= 16'h0500;
// mem[1781] <= 16'h0b00;
// mem[1782] <= 16'h0000;
// mem[1783] <= 16'h0700;
// mem[1784] <= 16'h0200;
// mem[1785] <= 16'h0500;
// mem[1786] <= 16'h0b00;
// mem[1787] <= 16'h0200;
// mem[1788] <= 16'hffff;
// mem[1789] <= 16'h0b00;
// mem[1790] <= 16'hfdff;
// mem[1791] <= 16'h0d00;
// mem[1792] <= 16'h0300;
// mem[1793] <= 16'h0400;
// mem[1794] <= 16'h0d00;
// mem[1795] <= 16'hf9ff;
// mem[1796] <= 16'h0d00;
// mem[1797] <= 16'hffff;
// mem[1798] <= 16'h0000;
// mem[1799] <= 16'h0300;
// mem[1800] <= 16'h0200;
// mem[1801] <= 16'h0600;
// mem[1802] <= 16'h0300;
// mem[1803] <= 16'h0200;
// mem[1804] <= 16'h0900;
// mem[1805] <= 16'h0300;
// mem[1806] <= 16'h0700;
// mem[1807] <= 16'hffff;
// mem[1808] <= 16'h0900;
// mem[1809] <= 16'hffff;
// mem[1810] <= 16'h0500;
// mem[1811] <= 16'h0900;
// mem[1812] <= 16'h0000;
// mem[1813] <= 16'h0700;
// mem[1814] <= 16'h0200;
// mem[1815] <= 16'h0500;
// mem[1816] <= 16'h0500;
// mem[1817] <= 16'h0000;
// mem[1818] <= 16'h0600;
// mem[1819] <= 16'hfbff;
// mem[1820] <= 16'h0200;
// mem[1821] <= 16'h0700;
// mem[1822] <= 16'h0200;
// mem[1823] <= 16'h0000;
// mem[1824] <= 16'h0200;
// mem[1825] <= 16'h0000;
// mem[1826] <= 16'hfdff;
// mem[1827] <= 16'h0b00;
// mem[1828] <= 16'h0000;
// mem[1829] <= 16'hfdff;
// mem[1830] <= 16'h0500;
// mem[1831] <= 16'h0500;
// mem[1832] <= 16'h0000;
// mem[1833] <= 16'h0500;
// mem[1834] <= 16'hfdff;
// mem[1835] <= 16'h0200;
// mem[1836] <= 16'h0700;
// mem[1837] <= 16'h0000;
// mem[1838] <= 16'h0900;
// mem[1839] <= 16'hfdff;
// mem[1840] <= 16'h0200;
// mem[1841] <= 16'h0700;
// mem[1842] <= 16'h0200;
// mem[1843] <= 16'hf9ff;
// mem[1844] <= 16'h0900;
// mem[1845] <= 16'h0300;
// mem[1846] <= 16'h0200;
// mem[1847] <= 16'h0200;
// mem[1848] <= 16'h0200;
// mem[1849] <= 16'h0200;
// mem[1850] <= 16'h0200;
// mem[1851] <= 16'h0700;
// mem[1852] <= 16'h0000;
// mem[1853] <= 16'h0200;
// mem[1854] <= 16'h0000;
// mem[1855] <= 16'hfdff;
// mem[1856] <= 16'h0200;
// mem[1857] <= 16'hf9ff;
// mem[1858] <= 16'h0600;
// mem[1859] <= 16'h0000;
// mem[1860] <= 16'hfdff;
// mem[1861] <= 16'h0000;
// mem[1862] <= 16'h0000;
// mem[1863] <= 16'h0200;
// mem[1864] <= 16'h0200;
// mem[1865] <= 16'hfdff;
// mem[1866] <= 16'hfdff;
// mem[1867] <= 16'h0700;
// mem[1868] <= 16'hffff;
// mem[1869] <= 16'h0200;
// mem[1870] <= 16'hfdff;
// mem[1871] <= 16'h0500;
// mem[1872] <= 16'hffff;
// mem[1873] <= 16'hf7ff;
// mem[1874] <= 16'h0000;
// mem[1875] <= 16'h0200;
// mem[1876] <= 16'h0000;
// mem[1877] <= 16'h0200;
// mem[1878] <= 16'h0000;
// mem[1879] <= 16'hf9ff;
// mem[1880] <= 16'h0500;
// mem[1881] <= 16'h0000;
// mem[1882] <= 16'h0000;
// mem[1883] <= 16'h0000;
// mem[1884] <= 16'hfbff;
// mem[1885] <= 16'h0300;
// mem[1886] <= 16'hffff;
// mem[1887] <= 16'hffff;
// mem[1888] <= 16'hffff;
// mem[1889] <= 16'h0000;
// mem[1890] <= 16'hfdff;
// mem[1891] <= 16'hfdff;
// mem[1892] <= 16'hf7ff;
// mem[1893] <= 16'h0800;
// mem[1894] <= 16'h0200;
// mem[1895] <= 16'hffff;
// mem[1896] <= 16'h0000;
// mem[1897] <= 16'h0200;
// mem[1898] <= 16'hf5ff;
// mem[1899] <= 16'h0200;
// mem[1900] <= 16'h0000;
// mem[1901] <= 16'h0000;
// mem[1902] <= 16'hf9ff;
// mem[1903] <= 16'h0200;
// mem[1904] <= 16'h0500;
// mem[1905] <= 16'hfbff;
// mem[1906] <= 16'hfdff;
// mem[1907] <= 16'hfbff;
// mem[1908] <= 16'hfbff;
// mem[1909] <= 16'hfdff;
// mem[1910] <= 16'hfbff;
// mem[1911] <= 16'h0500;
// mem[1912] <= 16'hf1ff;
// mem[1913] <= 16'h0500;
// mem[1914] <= 16'hfbff;
// mem[1915] <= 16'h0500;
// mem[1916] <= 16'hf7ff;
// mem[1917] <= 16'h0200;
// mem[1918] <= 16'hfdff;
// mem[1919] <= 16'hf9ff;
// mem[1920] <= 16'h0200;
// mem[1921] <= 16'h0200;
// mem[1922] <= 16'hf5ff;
// mem[1923] <= 16'hfdff;
// mem[1924] <= 16'hf7ff;
// mem[1925] <= 16'hffff;
// mem[1926] <= 16'h0200;
// mem[1927] <= 16'hf5ff;
// mem[1928] <= 16'h0300;
// mem[1929] <= 16'h0000;
// mem[1930] <= 16'hf5ff;
// mem[1931] <= 16'h0000;
// mem[1932] <= 16'h0000;
// mem[1933] <= 16'hfdff;
// mem[1934] <= 16'hfdff;
// mem[1935] <= 16'hfdff;
// mem[1936] <= 16'hfdff;
// mem[1937] <= 16'hfbff;
// mem[1938] <= 16'h0300;
// mem[1939] <= 16'hf7ff;
// mem[1940] <= 16'hf9ff;
// mem[1941] <= 16'h0300;
// mem[1942] <= 16'hfbff;
// mem[1943] <= 16'hfbff;
// mem[1944] <= 16'hffff;
// mem[1945] <= 16'hf7ff;
// mem[1946] <= 16'hffff;
// mem[1947] <= 16'hffff;
// mem[1948] <= 16'hf5ff;
// mem[1949] <= 16'hfdff;
// mem[1950] <= 16'h0200;
// mem[1951] <= 16'hffff;
// mem[1952] <= 16'hf5ff;
// mem[1953] <= 16'hffff;
// mem[1954] <= 16'hfbff;
// mem[1955] <= 16'hf9ff;
// mem[1956] <= 16'h0200;
// mem[1957] <= 16'hf9ff;
// mem[1958] <= 16'hfdff;
// mem[1959] <= 16'hf0ff;
// mem[1960] <= 16'hffff;
// mem[1961] <= 16'hfdff;
// mem[1962] <= 16'hf5ff;
// mem[1963] <= 16'h0300;
// mem[1964] <= 16'hf1ff;
// mem[1965] <= 16'h0000;
	end
end


endmodule // audio_loop
